`ifndef __PCSELECT_SV
`define __PCSELECT_SV

`ifdef VERILATOR
`include "include/common.sv"
`include "include/pipes.sv" 
`else

`endif 

module pcselect
import common::*;
import pipes::*;
(
    input u64 pcplus4,
    output u64 pc_selected,
    input u1 stall
);

    always_comb
    begin
        if(stall)
            pc_selected = pcplus4 - 4;
        else
            pc_selected = pcplus4;
    end

endmodule
`endif

